-----------------Laboratorio Digital-------------------------------------
-- Arquivo   : rom_angulos_141x24.vhd
-- Projeto   : Experiencia 6 - Sistema de Sonar
-------------------------------------------------------------------------
-- Descricao : 
--             memoria rom 16x24 (descricao comportamental)
--             conteudo com 16 posicoes angulares predefinidos
-------------------------------------------------------------------------
-- Revisoes  :
--     Data        Versao  Autor             Descricao
--     20/09/2019  1.0     Edson Midorikawa  criacao
--     01/10/2020  1.1     Edson Midorikawa  revisao
--     09/10/2021  1.2     Edson Midorikawa  revisao
--     24/09/2022  1.3     Edson Midorikawa  revisao
--     31/10/2022  2.0     Gabriel Zambelli  refatoraçao
-------------------------------------------------------------------------
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity rom_angulos_141x24 is
    port (
        endereco : in  std_logic_vector(9 downto 0);
        saida    : out std_logic_vector(23 downto 0)
    ); 
end entity;


architecture rom_arch of rom_angulos_141x24 is

    signal posicao_memoria: integer;

    type memoria_8x24 is array (integer range 0 to 140) of std_logic_vector(23 downto 0);

    constant tabela_angulos: memoria_8x24 := (
        x"303230", --     0 = 020  -- conteudo da ROM
        x"303231", --     1 = 021  -- angulos para o sonar
        x"303232", --     2 = 022  -- (valores em hexadecimal)
        x"303233", --     3 = 023
        x"303234", --     4 = 024
        x"303235", --     5 = 025
        x"303236", --     6 = 026
        x"303237", --     7 = 027
        x"303238", --     8 = 028
        x"303239", --     9 = 029
        x"303330", --    10 = 030
        x"303331", --    11 = 031
        x"303332", --    12 = 032
        x"303333", --    13 = 033
        x"303334", --    14 = 034
        x"303335", --    15 = 035
        x"303336", --    16 = 036
        x"303337", --    17 = 037
        x"303338", --    18 = 038
        x"303339", --    19 = 039
        x"303430", --    20 = 040
        x"303431", --    21 = 041
        x"303432", --    22 = 042
        x"303433", --    23 = 043
        x"303434", --    24 = 044
        x"303435", --    25 = 045
        x"303436", --    26 = 046
        x"303437", --    27 = 047
        x"303438", --    28 = 048
        x"303439", --    29 = 049
        x"303530", --    30 = 050
        x"303531", --    31 = 051
        x"303532", --    32 = 052
        x"303533", --    33 = 053
        x"303534", --    34 = 054
        x"303535", --    35 = 055
        x"303536", --    36 = 056
        x"303537", --    37 = 057
        x"303538", --    38 = 058
        x"303539", --    39 = 059
        x"303630", --    40 = 060
        x"303631", --    41 = 061
        x"303632", --    42 = 062
        x"303633", --    43 = 063
        x"303634", --    44 = 064
        x"303635", --    45 = 065
        x"303636", --    46 = 066
        x"303637", --    47 = 067
        x"303638", --    48 = 068
        x"303639", --    49 = 069
        x"303730", --    50 = 070
        x"303731", --    51 = 071
        x"303732", --    52 = 072
        x"303733", --    53 = 073
        x"303734", --    54 = 074
        x"303735", --    55 = 075
        x"303736", --    56 = 076
        x"303737", --    57 = 077
        x"303738", --    58 = 078
        x"303739", --    59 = 079
        x"303830", --    60 = 080
        x"303831", --    61 = 081
        x"303832", --    62 = 082
        x"303833", --    63 = 083
        x"303834", --    64 = 084
        x"303835", --    65 = 085
        x"303836", --    66 = 086
        x"303837", --    67 = 087
        x"303838", --    68 = 088
        x"303839", --    69 = 089
        x"303930", --    70 = 090
        x"303931", --    71 = 091
        x"303932", --    72 = 092
        x"303933", --    73 = 093
        x"303934", --    74 = 094
        x"303935", --    75 = 095
        x"303936", --    76 = 096
        x"303937", --    77 = 097
        x"303938", --    78 = 098
        x"303939", --    79 = 099
        x"313030", --    80 = 100
        x"313031", --    81 = 101
        x"313032", --    82 = 102
        x"313033", --    83 = 103
        x"313034", --    84 = 104
        x"313035", --    85 = 105
        x"313036", --    86 = 106
        x"313037", --    87 = 107
        x"313038", --    88 = 108
        x"313039", --    89 = 109
        x"313130", --    90 = 110
        x"313131", --    91 = 111
        x"313132", --    92 = 112
        x"313133", --    93 = 113
        x"313134", --    94 = 114
        x"313135", --    95 = 115
        x"313136", --    96 = 116
        x"313137", --    97 = 117
        x"313138", --    98 = 118
        x"313139", --    99 = 119
        x"313230", --   100 = 120
        x"313231", --   101 = 121
        x"313232", --   102 = 122
        x"313233", --   103 = 123
        x"313234", --   104 = 124
        x"313235", --   105 = 125
        x"313236", --   106 = 126
        x"313237", --   107 = 127
        x"313238", --   108 = 128
        x"313239", --   109 = 129
        x"313330", --   110 = 130
        x"313331", --   111 = 131
        x"313332", --   112 = 132
        x"313333", --   113 = 133
        x"313334", --   114 = 134
        x"313335", --   115 = 135
        x"313336", --   116 = 136
        x"313337", --   117 = 137
        x"313338", --   118 = 138
        x"313339", --   119 = 139
        x"313430", --   120 = 140
        x"313431", --   121 = 141
        x"313432", --   122 = 142
        x"313433", --   123 = 143
        x"313434", --   124 = 144
        x"313435", --   125 = 145
        x"313436", --   126 = 146
        x"313437", --   127 = 147
        x"313438", --   128 = 148
        x"313439", --   129 = 149
        x"313530", --   130 = 150
        x"313531", --   131 = 151
        x"313532", --   132 = 152
        x"313533", --   133 = 153
        x"313534", --   134 = 154
        x"313535", --   135 = 155
        x"313536", --   136 = 156
        x"313537", --   137 = 157
        x"313538", --   138 = 158
        x"313539", --   139 = 159
        x"313630"  --   140 = 160
    );

begin

    -- converte os 8 primeiros dígitos (2^8 = 256) para caber de 0 a 140
    posicao_memoria <= to_integer(unsigned(endereco(9 downto 2))) * 141 / 256;

    saida   <= tabela_angulos(posicao_memoria);

end architecture rom_arch;
